// SPDX-License-Identifier: CERN-OHL-P
// Copyright 2024 regymm
// Wrapped and configured pcie_7x for use with litepcie
`timescale 1ns / 1ps
`default_nettype wire

module pcie_s7 (
	// Tx
	output  [0:0] pci_exp_txn,
	output  [0:0] pci_exp_txp,
	// Rx
	input   [0:0] pci_exp_rxn,
	input   [0:0] pci_exp_rxp,
	input   pipe_mmcm_rst_n,
	output  pipe_mmcm_lock,
	// AXIS Common
	output                                     user_clk_out,
	output                                     user_reset_out,
	output                                     user_lnk_up,

	input                                      tx_cfg_gnt,
	input                                      rx_np_ok,
	input                                      rx_np_req,
	input                                      cfg_turnoff_ok,
	input                                      cfg_trn_pending,
	input                                      cfg_pm_halt_aspm_l0s,
	input                                      cfg_pm_halt_aspm_l1,
	input                                      cfg_pm_force_state_en,
	input    [1:0]                             cfg_pm_force_state,
	input    [63:0]                            cfg_dsn,
	input                                      cfg_pm_wake,
	// AXI TX
	input   [64-1:0]                           s_axis_tx_tdata,
	input                                      s_axis_tx_tvalid,
	output                                     s_axis_tx_tready,
	input   [8-1:0]                            s_axis_tx_tkeep,
	input                                      s_axis_tx_tlast,
	input   [3:0]                              s_axis_tx_tuser,
	// AXI RX
	output  [64-1:0]                           m_axis_rx_tdata,
	output                                     m_axis_rx_tvalid,
	input                                      m_axis_rx_tready,
	output  [8-1:0]                            m_axis_rx_tkeep,
	output                                     m_axis_rx_tlast,
	output  [21:0]                             m_axis_rx_tuser,
	// Configuration (CFG) Interface
	// EP and RP
	output                                     tx_err_drop,
	output                                     tx_cfg_req,
	output  [5:0]                              tx_buf_av,
	output   [15:0]                            cfg_status,
	output   [15:0]                            cfg_command,
	output   [15:0]                            cfg_dstatus,
	output   [15:0]                            cfg_dcommand,
	output   [15:0]                            cfg_lstatus,
	output   [15:0]                            cfg_lcommand,
	output   [15:0]                            cfg_dcommand2,
	output   [2:0]                             cfg_pcie_link_state,
	output                                     cfg_to_turnoff,
	output   [7:0]                             cfg_bus_number,
	output   [4:0]                             cfg_device_number,
	output   [2:0]                             cfg_function_number,

	output                                     cfg_pmcsr_pme_en,
	output   [1:0]                             cfg_pmcsr_powerstate,
	output                                     cfg_pmcsr_pme_status,
	output                                     cfg_received_func_lvl_rst,
	// EP Only
	input                                       cfg_interrupt,
	output                                      cfg_interrupt_rdy,
	input                                       cfg_interrupt_assert,
	input    [7:0]                              cfg_interrupt_di,
	output   [7:0]                              cfg_interrupt_do,
	output   [2:0]                              cfg_interrupt_mmenable,
	output                                      cfg_interrupt_msienable,
	output                                      cfg_interrupt_msixenable,
	output                                      cfg_interrupt_msixfm,
	input                                       cfg_interrupt_stat,
	input    [4:0]                              cfg_pciecap_interrupt_msgnum,

	input                                       sys_clk,
	input                                       sys_rst_n,
	output   [4:0]                              gt_reset_fsm,
	output   [5:0]                              pl_ltssm_state,

  // use external MMCM for litepcie
  input                                       pipe_pclk_in,
  input                                       pipe_dclk_in,
  input                                       pipe_oobclk_in,
  input                                       pipe_userclk1_in,
  input                                       pipe_userclk2_in,
  input                                       pipe_mmcm_lock_in,
  input                                       pipe_rxusrclk_in,
  input                                       pipe_rxoutclk_in,

  output                                      pipe_pclk_sel_out,
  output                                      pipe_txoutclk_out,

  // unused cfgs, if problem occur, connect it to block in pcie_7x
  input                                       cfg_aer_interrupt_msgnum,
  input                                       cfg_ds_bus_number,
  input                                       cfg_ds_device_number,
  input                                       cfg_ds_function_number,
  input                                       cfg_err_acs,
  input                                       cfg_err_aer_headerlog,
  input                                       cfg_err_atomic_egress_blocked,
  input                                       cfg_err_cor,
  input                                       cfg_err_cpl_abort,
  input                                       cfg_err_cpl_timeout,
  input                                       cfg_err_cpl_unexpect,
  input                                       cfg_err_ecrc,
  input                                       cfg_err_internal_cor,
  input                                       cfg_err_internal_uncor,
  input                                       cfg_err_locked,
  input                                       cfg_err_malformed,
  input                                       cfg_err_mc_blocked,
  input                                       cfg_err_norecovery,
  input                                       cfg_err_poisoned,
  input                                       cfg_err_posted,
  input                                       cfg_err_tlp_cpl_header,
  input                                       cfg_err_ur,
  input                                       cfg_mgmt_byte_en,
  input                                       cfg_mgmt_di,
  input                                       cfg_mgmt_dwaddr,
  input                                       cfg_mgmt_rd_en,
  input                                       cfg_mgmt_wr_en,
  input                                       cfg_mgmt_wr_readonly,
  input                                       cfg_mgmt_wr_rw1c_as_rw,
  input                                       cfg_pm_send_pme_to,
  input                                       fc_sel,
  input                                       pcie_drp_addr,
  input                                       pcie_drp_clk,
  input                                       pcie_drp_di,
  input                                       pcie_drp_en,
  input                                       pcie_drp_we,
  input                                       pl_directed_link_auton,
  input                                       pl_directed_link_change,
  input                                       pl_directed_link_speed,
  input                                       pl_directed_link_width,
  input                                       pl_downstream_deemph_source,
  input                                       pl_transmit_hot_rst,
  input                                       pl_upstream_prefer_deemph,

  output                                      cfg_aer_ecrc_check_en,
  output                                      cfg_aer_ecrc_gen_en,
  output                                      cfg_aer_rooterr_corr_err_received,
  output                                      cfg_aer_rooterr_corr_err_reporting_en,
  output                                      cfg_aer_rooterr_fatal_err_received,
  output                                      cfg_aer_rooterr_fatal_err_reporting_en,
  output                                      cfg_aer_rooterr_non_fatal_err_received,
  output                                      cfg_aer_rooterr_non_fatal_err_reporting_en,
  output                                      cfg_bridge_serr_en,
  output                                      cfg_err_aer_headerlog_set,
  output                                      cfg_err_cpl_rdy,
  output                                      cfg_mgmt_do,
  output                                      cfg_mgmt_rd_wr_done,
  output                                      cfg_msg_data,
  output                                      cfg_msg_received,
  output                                      cfg_msg_received_assert_int_a,
  output                                      cfg_msg_received_assert_int_b,
  output                                      cfg_msg_received_assert_int_c,
  output                                      cfg_msg_received_assert_int_d,
  output                                      cfg_msg_received_deassert_int_a,
  output                                      cfg_msg_received_deassert_int_b,
  output                                      cfg_msg_received_deassert_int_c,
  output                                      cfg_msg_received_deassert_int_d,
  output                                      cfg_msg_received_err_cor,
  output                                      cfg_msg_received_err_fatal,
  output                                      cfg_msg_received_err_non_fatal,
  output                                      cfg_msg_received_pm_as_nak,
  output                                      cfg_msg_received_pm_pme,
  output                                      cfg_msg_received_pme_to_ack,
  output                                      cfg_msg_received_setslotpowerlimit,
  output                                      cfg_root_control_pme_int_en,
  output                                      cfg_root_control_syserr_corr_err_en,
  output                                      cfg_root_control_syserr_fatal_err_en,
  output                                      cfg_root_control_syserr_non_fatal_err_en,
  output                                      cfg_slot_control_electromech_il_ctl_pulse,
  output                                      cfg_vc_tcvc_map,
  output                                      fc_cpld,
  output                                      fc_cplh,
  output                                      fc_npd,
  output                                      fc_nph,
  output                                      fc_pd,
  output                                      fc_ph,
  output                                      pcie_drp_do,
  output                                      pcie_drp_rdy,
  output                                      pipe_gen3_out,
  output                                      pipe_rxoutclk_out,
  output                                      pl_directed_change_done,
  output                                      pl_initial_link_width,
  output                                      pl_lane_reversal_mode,
  output                                      pl_link_gen2_cap,
  output                                      pl_link_partner_gen2_supported,
  output                                      pl_link_upcfg_cap,
  output                                      pl_phy_lnk_up,
  output                                      pl_received_hot_rst,
  output                                      pl_rx_pm_state,
  output                                      pl_sel_lnk_rate,
  output                                      pl_sel_lnk_width,
  output                                      pl_tx_pm_state,
  output                                      user_app_rdy
);

pcie_7x #(
  .EXTERNAL_MMCM("TRUE"),
  .BAR0(32'hFC000000),
  .USER_CLK_FREQ(2)
) pcie_7x_litepcie_inst (
  .pci_exp_txn(pci_exp_txn),
  .pci_exp_txp(pci_exp_txp),
  .pci_exp_rxn(pci_exp_rxn),
  .pci_exp_rxp(pci_exp_rxp),
  .pipe_mmcm_rst_n(pipe_mmcm_rst_n),
  .pipe_mmcm_lock(pipe_mmcm_lock),
  
  .user_clk_out(user_clk_out),
  .user_reset_out(user_reset_out),
  .user_lnk_up(user_lnk_up),

  .tx_cfg_gnt(tx_cfg_gnt),
  .rx_np_ok(rx_np_ok),
  .rx_np_req(rx_np_req),
  .cfg_turnoff_ok(cfg_turnoff_ok),
  .cfg_trn_pending(cfg_trn_pending),
  .cfg_pm_halt_aspm_l0s(cfg_pm_halt_aspm_l0s),
  .cfg_pm_halt_aspm_l1(cfg_pm_halt_aspm_l1),
  .cfg_pm_force_state_en(cfg_pm_force_state_en),
  .cfg_pm_force_state(cfg_pm_force_state),
  .cfg_dsn(cfg_dsn),
  .cfg_pm_wake(cfg_pm_wake),

  .s_axis_tx_tdata(s_axis_tx_tdata),
  .s_axis_tx_tvalid(s_axis_tx_tvalid),
  .s_axis_tx_tready(s_axis_tx_tready),
  .s_axis_tx_tkeep(s_axis_tx_tkeep),
  .s_axis_tx_tlast(s_axis_tx_tlast),
  .s_axis_tx_tuser(s_axis_tx_tuser),

  .m_axis_rx_tdata(m_axis_rx_tdata),
  .m_axis_rx_tvalid(m_axis_rx_tvalid),
  .m_axis_rx_tready(m_axis_rx_tready),
  .m_axis_rx_tkeep(m_axis_rx_tkeep),
  .m_axis_rx_tlast(m_axis_rx_tlast),
  .m_axis_rx_tuser(m_axis_rx_tuser),

  .tx_err_drop(tx_err_drop),
  .tx_cfg_req(tx_cfg_req),
  .tx_buf_av(tx_buf_av),
  .cfg_status(cfg_status),
  .cfg_command(cfg_command),
  .cfg_dstatus(cfg_dstatus),
  .cfg_dcommand(cfg_dcommand),
  .cfg_lstatus(cfg_lstatus),
  .cfg_lcommand(cfg_lcommand),
  .cfg_dcommand2(cfg_dcommand2),
  .cfg_pcie_link_state(cfg_pcie_link_state),
  .cfg_to_turnoff(cfg_to_turnoff),
  .cfg_bus_number(cfg_bus_number),
  .cfg_device_number(cfg_device_number),
  .cfg_function_number(cfg_function_number),
  .cfg_pmcsr_pme_en(cfg_pmcsr_pme_en),
  .cfg_pmcsr_powerstate(cfg_pmcsr_powerstate),
  .cfg_pmcsr_pme_status(cfg_pmcsr_pme_status),
  .cfg_received_func_lvl_rst(cfg_received_func_lvl_rst),
  .cfg_interrupt(cfg_interrupt),
  .cfg_interrupt_rdy(cfg_interrupt_rdy),
  .cfg_interrupt_assert(cfg_interrupt_assert),
  .cfg_interrupt_di(cfg_interrupt_di),
  .cfg_interrupt_do(cfg_interrupt_do),
  .cfg_interrupt_mmenable(cfg_interrupt_mmenable),
  .cfg_interrupt_msienable(cfg_interrupt_msienable),
  .cfg_interrupt_msixenable(cfg_interrupt_msixenable),
  .cfg_interrupt_msixfm(cfg_interrupt_msixfm),
  .cfg_interrupt_stat(cfg_interrupt_stat),
  .cfg_pciecap_interrupt_msgnum(cfg_pciecap_interrupt_msgnum),

  .sys_clk(sys_clk),
  .sys_rst_n(sys_rst_n),
  .gt_reset_fsm(),
  .pl_ltssm_state(pl_ltssm_state),

  .pipe_pclk_in(pipe_pclk_in),
  .pipe_dclk_in(pipe_dclk_in),
  .pipe_oobclk_in(pipe_oobclk_in),
  .pipe_userclk1_in(pipe_userclk1_in),
  .pipe_userclk2_in(pipe_userclk2_in),
  .pipe_mmcm_lock_in(pipe_mmcm_lock_in),
  .pipe_rxusrclk_in(pipe_rxusrclk_in),
  .pipe_rxoutclk_in(pipe_rxoutclk_in),
  .pipe_pclk_sel_out(pipe_pclk_sel_out),
  .pipe_txoutclk_out(pipe_txoutclk_out)
);

endmodule
